module dmem_sel (
    input [31:0] addr,
    input [31:0] din,
    input [2:0] funct3,
	input pc30,
    output [31:0] dout,
    output [11:0] bios_addrb,
    input [31:0] bios_doutb,
    output [13:0] dmem_addra,
    output [31:0] dmem_dina,
    output [3:0] dmem_wea,
    input [31:0] dmem_douta,
    output [13:0] imem_addra,
    output [31:0] imem_dina,
    output [3:0] imem_wea
);

    assign bios_addrb = addr[11:0];
    assign dmem_addra = addr[13:0];
    assign imem_addra = addr[13:0];
    assign dmem_dina = din;
    assign imem_dina = din;
    
	
    reg [3:0] wea;
    
    always @ (*) begin
        case (funct3)
            FNC_SB:
                case (addr[1:0])
                    2'b00:
                        wea = 4'b0001;
                    2'b01:
                        wea = 4'b0010;
                    2'b10:
                        wea = 4'b0100;
                    2'b11:
                        wea = 4'b1000;
                endcase
            FNC_SH:
                case (addr[1])
                    2'b0:
                        wea = 4'b0011;
                    2'b1:
                        wea = 4'b1100;
                endcase
            FNC_SW:
                wea = 4'b1111;
            default:
                wea = 4'b0000;
        endcase
    end

    assign dmem_wea = addr[28] == 1'b1 ? wea : 4'b0000;
    assign imem_wea = addr[29] == 1'b1 && pc30 == 1'b1 ? wea : 4'b0000;
    assign dout = addr[31:28] == 4'b0100 ? bios_doutb : dmem_douta;

endmodule